`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 17.03.2022 19:37:32
// Design Name: 
// Module Name: Output_layer
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Output_layer(
    input wire ,
    input wire [15:0] V,
    output wire [15:0] y
    );

reg [7:0] W_out [0:49];

    
    
endmodule
