`timescale 1ns / 1ps


module Output_layer(
    input wire ,
    input wire [15:0] V,
    output wire [15:0] y
    );

reg [7:0] W_out [0:49];

    
    
endmodule
